/* 
 * mac_ctrl.sv
 * Francesco Conti <fconti@iis.ee.ethz.ch>
 *
 * Copyright (C) 2018 ETH Zurich, University of Bologna
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 */

import mac_package::*;
import hwpe_ctrl_package::*;

module mac_ctrl
#(
  parameter int unsigned N_CORES         = 2,
  parameter int unsigned N_CONTEXT       = 2,
  parameter int unsigned N_IO_REGS       = 17, 
  parameter int unsigned ID              = 10,
  parameter int unsigned UCODE_HARDWIRED = 0 //if this is 1, then ucode_flat will be equal to the code generated by ucode_compile.py 
)
(
  // global signals
  input  logic                                  clk_i,
  input  logic                                  rst_ni,
  input  logic                                  test_mode_i,
  output logic                                  clear_o,
  // events
  output logic [N_CORES-1:0][REGFILE_N_EVT-1:0] evt_o, //parameter REGFILE_N_EVT defined in hwpe_ctrl_package
  // ctrl & flags
  output ctrl_streamer_t                        ctrl_streamer_o,
  input  flags_streamer_t                       flags_streamer_i,
  output ctrl_engine_t                          ctrl_engine_o,
  input  flags_engine_t                         flags_engine_i,
  // periph slave port
  hwpe_ctrl_intf_periph.slave                   periph
);

  ctrl_slave_t   slave_ctrl;
  flags_slave_t  slave_flags;
  ctrl_regfile_t reg_file; //important to program microcontroller work as it should

  logic unsigned [31:0] static_reg_nb_if;
  logic unsigned [31:0] static_reg_nb_of;
  //logic unsigned [31:0] static_reg_ow_x_nof;
  logic unsigned [31:0] static_reg_iw_x_nif;
  logic unsigned [31:0] static_reg_nfa;
  logic unsigned [31:0] static_reg_nwa;
  logic unsigned [31:0] static_reg_zero;
  logic unsigned [31:0] static_reg_nfw;
  logic unsigned [31:0] static_reg_loop1_loop0;
  logic unsigned [31:0] static_reg_loop3_loop2;
  logic unsigned [31:0] static_reg_loop5_loop4;
  logic unsigned [31:0] static_reg_cnt_prog1;
  logic unsigned [31:0] static_reg_cnt_prog2;
  logic unsigned [31:0] static_reg_iter_len_wei_out;
  logic unsigned [31:0] static_reg_par_sel;

  logic [223:0]  ucode_flat;
  ucode_t ucode;
  ctrl_ucode_t   ucode_ctrl;
  flags_ucode_t  ucode_flags;
  logic [11:0][31:0] ucode_registers_read; //of course, you have 12 RO registers with size 32 bits, here just use the ones you need

  ctrl_fsm_t fsm_ctrl;

  /* Peripheral slave & register file */
  hwpe_ctrl_slave #(
    .N_CORES        ( N_CORES               ),
    .N_CONTEXT      ( N_CONTEXT             ),
    .N_IO_REGS      ( N_IO_REGS             ),
    .N_GENERIC_REGS ( (1-UCODE_HARDWIRED)*8 ),
    .ID_WIDTH       ( ID                    )
  ) i_slave (
    .clk_i    ( clk_i       ),
    .rst_ni   ( rst_ni      ),
    .clear_o  ( clear_o     ),
    .cfg      ( periph      ),
    .ctrl_i   ( slave_ctrl  ),
    .flags_o  ( slave_flags ),
    .reg_file ( reg_file    )
  );
  assign evt_o = slave_flags.evt;

  /* Direct register file mappings */
  assign static_reg_nb_if      		= reg_file.hwpe_params[MAC_REG_NIF]; 
  assign static_reg_nb_of    		= reg_file.hwpe_params[MAC_REG_NOF];
  //assign static_reg_ow_x_nof   	= reg_file.hwpe_params[MAC_REG_OW_X_NOF];
  assign static_reg_iw_x_nif   		= reg_file.hwpe_params[MAC_REG_IW_X_NIF];
  assign static_reg_nfa     		= reg_file.hwpe_params[MAC_REG_NFA];
  assign static_reg_nwa  		= reg_file.hwpe_params[MAC_REG_NWA];
  assign static_reg_zero		= reg_file.hwpe_params[MAC_REG_ZERO];
  assign static_reg_nfw			= reg_file.hwpe_params[MAC_REG_NFW];
  //to the following loops a +1 is added because this allows to extend the counting range
  //during accelerator programming take this into account when loading up the register file 
  assign static_reg_loop1_loop0		= reg_file.hwpe_params[MAC_REG_LOOP1_LOOP0]+32'h00010001; //correggi spacchetta e ricompatta
  assign static_reg_loop3_loop2		= reg_file.hwpe_params[MAC_REG_LOOP3_LOOP2]+32'h00010001;
  assign static_reg_loop5_loop4		= reg_file.hwpe_params[MAC_REG_LOOP5_LOOP4]+32'h00010001;
  //these are needed by low level fsm
  assign static_reg_cnt_prog1  		= reg_file.hwpe_params[MAC_REG_CNT_PROG1];
  assign static_reg_cnt_prog2  		= reg_file.hwpe_params[MAC_REG_CNT_PROG2];	
  //these are needed by high level fsm
  assign static_reg_iter_len_wei_out 	= reg_file.hwpe_params[MAC_REG_ITER_LEN_WEI_OUT];
  assign static_reg_par_sel= reg_file.hwpe_params[MAC_REG_PAR_SEL]; 
  
  /* Microcode processor */
  generate
    if(UCODE_HARDWIRED) begin
      // equivalent to the microcode in ucode/code.yml (copy code generated by ucode_compile.py: first 176 are tail, rest is head)
      assign ucode_flat = 224'h5a432b2112020000000046788c02a3244504712205c278490121440b;
    end
    else begin
      // the microcode is stored in registers independent of context (job): in the testbench, during start-up you will have to 
	  // store the equivalent to the microcode in ucode/code.yml generated by ucode_compile.py in groups of 8 each (each generic reg is
	  //32 bit wide!)
      assign ucode_flat = reg_file.generic_params[6:0];
    end
  endgenerate
  
  assign ucode = { 
    // loops & bytecode
    ucode_flat,
    // loop ranges from outermost to innermost
    static_reg_loop5_loop4[27:16],
    static_reg_loop5_loop4[11:0],
    static_reg_loop3_loop2[27:16],
    static_reg_loop3_loop2[11:0],
    static_reg_loop1_loop0[27:16],
    static_reg_loop1_loop0[11:0]
  };
  
  //the following assignments are to program the programmable counter in the low level control inside the engine mac_engine.sv
  //the fileds into the two registers where values are saved are taken "randomly" but leaving enough space for the "parametric fields"
  assign ctrl_engine_o.max_val_in_vol 	              = static_reg_cnt_prog1[$clog2(MNV)-1:0];	 	 //no more than 26 bits
  assign ctrl_engine_o.max_val_cnt_relu_and_fil_group = static_reg_cnt_prog1[28:26];
  assign ctrl_engine_o.max_val_cnt_out 		      = static_reg_cnt_prog1[31:29];				
  assign ctrl_engine_o.max_val_cnt_done		      = static_reg_cnt_prog2[$clog2(MNO)-1:0]; 		 //no more than 25 bits
  assign ctrl_engine_o.max_val_cnt_quant 	      = static_reg_cnt_prog2[$clog2(Pa*Pw)-1+25:25]; //no more than 7 bits
  assign ctrl_engine_o.par_sel_Pa               = static_reg_par_sel[2]; //activations parallelism selection
  assign ctrl_engine_o.par_sel_Pw               = static_reg_par_sel[1:0]; //weights parallelism selection
 
  //start signal sent to the low level FSM
  //assign ctrl_engine_o.start = slave_flags.start;
 
  //the following assignments are for the RO registers in the ucontroller's RF
  assign ucode_registers_read[MAC_UCODE_MNEM_NIF]     	= static_reg_nb_if;
  assign ucode_registers_read[MAC_UCODE_MNEM_NOF] 	= static_reg_nb_of;
  //assign ucode_registers_read[MAC_UCODE_MNEM_OW_X_NOF]  = static_reg_ow_x_nof;
  assign ucode_registers_read[MAC_UCODE_MNEM_IW_X_NIF]  = static_reg_iw_x_nif;
  assign ucode_registers_read[MAC_UCODE_MNEM_NFA]  	= static_reg_nfa;
  assign ucode_registers_read[MAC_UCODE_MNEM_NWA]  	= static_reg_nwa;
  assign ucode_registers_read[MAC_UCODE_MNEM_ZERO]  	= static_reg_zero;
  assign ucode_registers_read[MAC_UCODE_MNEM_NFW] 	= static_reg_nfw;
  //the remaining registers are just filled with 0
  assign ucode_registers_read[11:7] = '0;
    
  
  hwpe_ctrl_ucode #(
    .NB_LOOPS  ( 6  ), //this is th enumber of loops to be supported (modified to 6)
    .NB_REG    ( 4  ), //this is the number of R/W registers
    .NB_RO_REG ( 12 )  //this is the number of read only registers
  ) i_ucode (
    .clk_i            ( clk_i                ),
    .rst_ni           ( rst_ni               ),
    .test_mode_i      ( test_mode_i          ),
    .clear_i          ( clear_o              ),
    .ctrl_i           ( ucode_ctrl           ),
    .flags_o          ( ucode_flags          ),
    .ucode_i          ( ucode                ),
    .registers_read_i ( ucode_registers_read )
  );

  /* Main FSM */
  mac_fsm i_fsm (
    .clk_i            ( clk_i              ),
    .rst_ni           ( rst_ni             ),
    .test_mode_i      ( test_mode_i        ),
    .clear_i          ( clear_o            ),
    .ctrl_streamer_o  ( ctrl_streamer_o    ),
    .flags_streamer_i ( flags_streamer_i   ),
    //.ctrl_engine_o    ( ctrl_engine_o      ), //not generated by top FSM
    .flags_engine_i   ( flags_engine_i     ),
    .ctrl_ucode_o     ( ucode_ctrl         ),
    .flags_ucode_i    ( ucode_flags        ),
    .ctrl_slave_o     ( slave_ctrl         ),
    .flags_slave_i    ( slave_flags        ),
    .reg_file_i       ( reg_file           ),
    .ctrl_i           ( fsm_ctrl           )
  );
  
  //the following must be changed according to your FSM: these are the lengths sent to top FSM to change the transaction size
  //and the line length of the generated addresses: these are used as number of 128 bits packets that will be fetched from or written to memory
  always_comb
  begin
    fsm_ctrl.len_wei        = static_reg_iter_len_wei_out[$clog2(MAC_CNT_LEN):0];     //(4*8*numfil/64) 
    fsm_ctrl.len_out        = static_reg_iter_len_wei_out[$clog2(MAC_CNT_LEN)+16:16]; //(4*num filtri/64)
  end

endmodule // mac_ctrl
