`timescale 1ns/1ns
//06/03/2019 this module is the top containing Data path and control unit
//this has been used just for synthesis purposes

import basic_package::*;
						 
module top 
	  #(parameter Pa = 8, 
		parameter Pw = 4,
		parameter M = 16,
		parameter BW = 128,
		parameter MNO = 288, 
		parameter MNV = 224*224)
	(	input clk,
		input rst_n,
		input core_stall_n,
		input [$clog2(MNO)-1:0] max_val_cnt_done,
		input [$clog2(Pa*Pw)-1:0] max_val_cnt_quant,
		input [2:0] max_val_cnt_out, max_val_cnt_relu, max_val_fil_group,
		input [$clog2(MNV)-1:0] max_val_in_vol,
		
		input [BW-1:0] in_data, 
		output [BW-1:0] out_data);	
	
	
	wire  w_en_mod_a, s_en_mod_a, act_load, w_en_a, w_en_w, w_en_br, MSB_a, w_and_s_ac1, cl_en_ac1, MSB_w, 
	      w_en_neg, valid_ac2, cl_en_ac2, valid_ac3, wb, cl_en_gen, s_en_ac3, cl_en_ac3; 
	wire [1:0] sel_mux_ac, sel_mux_out, sel_mux_relu;
	wire [7:0] wei_in_SMAC_reg_enables;

	CTRL_unit #(.Pa(Pa), .Pw(Pw), .MNO(MNO), .MNV(MNV)) controllo (
		.clk(clk), 
		.rst_n(rst_n), 
		.core_stall_n(core_stall_n),
		.max_val_cnt_done(max_val_cnt_done),
		.max_val_cnt_quant(max_val_cnt_quant),
		.max_val_cnt_out(max_val_cnt_out), 
		.max_val_cnt_relu(max_val_cnt_relu), 
		.max_val_fil_group(max_val_fil_group),
		.max_val_in_vol(max_val_in_vol),
		.act_load(act_load), 
		.w_en_mod_a(w_en_mod_a), 
		.s_en_mod_a(s_en_mod_a), 
		.w_en_a(w_en_a), 
		.w_en_w(w_en_w), 
		.w_en_br(w_en_br), 
		.MSB_a(MSB_a), 
		.w_and_s_ac1(w_and_s_ac1), 
		.cl_en_ac1(cl_en_ac1), 
		.MSB_w(MSB_w),
		.w_en_neg(w_en_neg), 
		.valid_ac2(valid_ac2), 
		.cl_en_ac2(cl_en_ac2), 
		.valid_ac3(valid_ac3), 
		.cl_en_ac3(cl_en_ac3), 
		.wb(wb), 
		.cl_en_gen(cl_en_gen), 
		.s_en_ac3(s_en_ac3),
		.sel_mux_out(sel_mux_out), 
		.sel_mux_relu(sel_mux_relu), 
		.sel_mux_ac(sel_mux_ac),
		.wei_in_SMAC_reg_enables(wei_in_SMAC_reg_enables)//,
		//temporary
		//.out_state(out_state)
	);
	
	Data_Path_1x64 #(.M(M), .Pa(Pa), .Pw(Pw), .MNO(MNO), .BW(BW)) Data_Path (
		.clk(clk), 
		.rst_n(rst_n),  
		.w_en_mod_a(w_en_mod_a), 
		.s_en_mod_a(s_en_mod_a), 
		.act_load(act_load),
		.cl_en_gen(cl_en_gen), 
		.w_en_a(w_en_a), 
		.w_en_w(w_en_w), 
		.w_en_br(w_en_br), 
		.MSB_a(MSB_a),
		.w_and_s_ac1(w_and_s_ac1), 
		.cl_en_ac1(cl_en_ac1), 
		.MSB_w(MSB_w), 
		.w_en_neg(w_en_neg), 
		.valid_ac2(valid_ac2), 
		.cl_en_ac2(cl_en_ac2),
		.valid_ac3(valid_ac3),  
		.wb(wb), 
		.s_en_ac3(s_en_ac3), 
		.cl_en_ac3(cl_en_ac3),
		.sel_mux_ac(sel_mux_ac),
		.sel_mux_relu(sel_mux_relu),
		.sel_mux_out(sel_mux_out), 
		.wei_in_SMAC_reg_enables(wei_in_SMAC_reg_enables),
		.in_data(in_data),
		.out_data(out_data)//,
		//TEMPORARY
		//.br_to_ac1_view(br_to_ac1_view),
		//.ac1_to_neg_view(ac1_to_neg_view),
		//.neg_to_ac2_view(neg_to_ac2_view),
		//.ac2_to_ac3_view(ac2_to_ac3_view),
		//.ac3_to_q_view(ac3_to_q_view)
	); 
	
	
	
endmodule
			
			